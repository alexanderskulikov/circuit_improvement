8 25 4
x0 x1 x2 x3 x4 x5 x6 x7
z0 x0 x1 0110
z1 x2 x3 0110
z2 x4 x5 0110
z3 x6 x7 0110
z4 z0 x0 0111
z5 z4 z0 0110
z6 x2 z0 0110
z7 z0 z1 0110
z8 z6 z1 0010
z9 z4 z8 0110
z10 x4 z7 0110
z11 z2 z10 0111
z12 z2 z7 0110
z13 z11 z12 0110
z14 x6 z12 0110
z15 z12 z3 0110
z16 z14 z3 0010
z17 z11 z16 0110
z18 z9 z5 0111
z19 z18 z9 0110
z20 z13 z9 0110
z21 z9 z17 0110
z22 z20 z17 0010
z23 z18 z22 0110
z24 z19 z23 0010
z15 z21 z23 z24