9 27 4
x1 x2 x3 x4 x5 x6 x7 x8 x9
z0 x1 x2 0110
z1 x2 x3 0110
z2 z0 z1 0111
z3 z0 x3 0110
z4 z2 z3 0110
z5 x4 z3 0110
z6 x4 x5 0110
z7 z5 z6 0010
z8 z3 z6 0110
z9 z2 z7 0110
z10 z4 z9 0010
z11 z8 x6 0110
z12 x6 x7 0110
z13 z11 z12 0111
z14 z11 x7 0110
z15 z13 z14 0110
z16 x8 z14 0110
z17 x8 x9 0110
z18 z16 z17 0010
z19 z14 z17 0110
z20 z13 z18 0110
z21 z15 z20 0010
z22 z9 z20 0110
z23 z9 z20 0001
z24 z10 z21 0110
z25 z23 z24 0110
z26 z10 z21 0001
z19 z22 z25 z26