5 11 1
x1 x2 x3 x4 x5
z1 x4 x5 0110
z2 x2 x3 1001
z4 z1 z2 1011
z7 x5 x3 1101
z8 x5 x4 1000
z10 x2 b6 0111
z11 x1 z10 1000
a9 z11 b8 1000
b6 z7 z8 0010
b7 x1 b6 1110
b8 z4 b7 0100
a9