15 51 4
x1 x2 x3 x4 x5 x6 x7 x8 x9 x10 x11 x12 x13 x14 x15 
2548 x5 x4 1001
1724 x12 4091 1001
4091 x10 4201 0110
4201 x11 5407 0110
5407 x9 5357 0110
5357 x8 5356 0110
5356 3591 x7 0110
4528 5297 3922 1001
5297 x2 x3 0110
3922 x1 2548 0110
457 x11 x10 0110
2056 5137 4806 0111
5137 5191 5301 1001
4806 5300 5027 0110
5191 5298 5355 0110
5301 5132 5300 1001
5300 5355 5299 1110
5027 5025 5409 1000
5298 5187 5296 0110
5355 5353 5354 1001
5132 4916 4142 1110
5299 4310 5298 1001
5025 5465 5191 0110
5409 5407 5408 0110
5187 5297 x1 0001
5296 x2 x3 0001
5353 3591 5352 0111
5354 4529 2548 0100
4916 5463 5465 1110
4142 5463 5246 0111
4310 5353 4528 1001
5246 5243 5244 1001
5243 1724 5242 0100
5244 1724 x13 0110
3652 457 4201 1000
4532 4527 5357 1110
4527 x8 x9 1001
3591 x6 4528 1001
5352 x7 x6 0110
4529 x4 4528 0110
2492 x14 x15 0110
5242 x12 x13 1001
3981 2056 4805 0110
4805 5301 5027 0110
5408 5191 4532 1001
5461 5244 x15 1001
5462 2492 5461 1000
5463 5243 5462 1001
5464 2492 5244 0110
5465 3652 5408 1001
5466 5463 5465 1001
5464 5466 4805 3981 