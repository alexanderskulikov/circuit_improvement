4 10 2
0 1 2 3
s4 0 1 1011
s5 1 2 0110
s6 s4 s5 1101
s7 2 s6 0010
s8 s5 s7 0110
s9 0 s8 0110
s10 s6 s9 1101
s11 3 s10 1001
s12 s6 s11 1110
s13 s9 s12 1011
s11 s13 