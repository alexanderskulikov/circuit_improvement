4 5 1
a b c d
e4 b d 0110
e5 d c 0110
e6 e4 e5 0100
e7 c e6 0110
e8 a e7 0111
e8