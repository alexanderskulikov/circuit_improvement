4 7 1
x1 x2 x3 x4
c5 x2 x1 0110
b6 d6 c8 0010
c8 x4 d5 0100
d3 c5 x2 1011
d4 c5 x3 1110
d5 x3 d3 1101
d6 d3 d4 0110
b6