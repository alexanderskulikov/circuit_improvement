6 13 1
x1 x2 x3 x4 x5 x6
z0 x1 x2 1001
z1 x1 x2 1000
z2 z1 x3 1001
z3 z0 z2 1001
z4 z1 z3 0100
z5 x4 z2 1001
z6 z5 z4 0111
z7 x5 z6 0110
z8 z7 z4 0110
z9 z8 x4 0110
z10 z9 z6 0001
z11 x6 z7 1001
z12 z10 z11 1000
z12