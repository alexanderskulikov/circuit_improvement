7 20 3
x1 x2 x3 x4 x5 x6 x7 
z0 x1 x2 0110
z1 x2 x3 0110
z2 z0 z1 0111
z3 z0 x3 0110
z4 z2 z3 0110
z5 z3 x4 0110
z6 x4 x5 0110
z7 z5 z6 0111
z8 z5 x5 0110
z9 z7 z8 0110
z10 z8 x6 0110
z11 x6 x7 0110
z12 z10 z11 0111
z13 z10 x7 0110
z14 z12 z13 0110
z15 z4 z9 0110
z16 z9 z14 0110
z17 z15 z16 0111
z18 z15 z14 0110
z19 z17 z18 0110
z13 z18 z19 