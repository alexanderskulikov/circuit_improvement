4 6 1
x1 x2 x3 x4 
z0 x2 x1 0010
z1 x4 x3 0001
z2 z0 z1 0111
z3 x4 x3 0111
z4 x1 z3 0100
z5 z2 z4 0110
z5 