8 18 2
x1 x2 x3 x4 x5 x6 x7 x8 
z0 x3 x2 1001
z1 z0 x1 0111
z2 z1 x4 0110
z3 z2 x1 0110
z4 z3 x3 0110
z5 z4 z1 0001
z6 z5 x5 1001
z7 z2 z6 1001
z8 z5 z7 0100
z9 x6 z6 1001
z10 z9 z8 0111
z11 z10 x7 0110
z12 z11 z8 0110
z13 z12 x6 0110
z14 z13 z10 0001
z15 z14 x8 1001
z16 z11 z15 1001
z17 z14 z16 0100
z17 z15 