16 83 16
x1 x2 x3 x4 x5 x6 x7 x8 x9 x10 x11 x12 x13 x14 x15 x16
z0 x4 x5 0110
z1 x6 x7 0110
z2 x8 x9 0110
z3 x10 x11 0110
z4 x12 x13 0110
z5 x14 x15 0110
z6 x1 x2 0110
z7 z6 x3 0110
z8 x1 x2 0001
z9 z6 x3 0001
z10 z8 z9 0110
z11 x4 z7 0110
z12 z0 z11 0111
z13 z0 z7 0110
z14 z12 z13 0110
z15 x6 z13 0110
z16 z13 z1 0110
z17 z15 z1 0010
z18 z12 z17 0110
z19 x8 z16 0110
z20 z2 z19 0111
z21 z2 z16 0110
z22 z20 z21 0110
z23 x10 z21 0110
z24 z21 z3 0110
z25 z23 z3 0010
z26 z20 z25 0110
z27 x12 z24 0110
z28 z4 z27 0111
z29 z4 z24 0110
z30 z28 z29 0110
z31 x14 z29 0110
z32 z29 z5 0110
z33 z31 z5 0010
z34 z28 z33 0110
z35 z14 z10 0110
z36 z18 z35 0111
z37 z18 z10 0110
z38 z36 z37 0110
z39 z22 z37 0110
z40 z37 z26 0110
z41 z39 z26 0010
z42 z36 z41 0110
z43 z40 z34 0110
z44 z30 z34 0010
z45 z40 z34 0001
z46 z44 z45 0110
z47 z46 z42 0110
z48 z38 z42 0010
z49 z46 z42 0001
z50 z48 z49 0110
z51 z32 x16 0110
z52 z32 x16 0001
z53 z43 z52 0110
z54 z43 z52 0001
z55 z47 z54 0110
z56 z47 z54 0001
z57 z50 z56 0110
a6 z53 z55 0001
a7 z55 vinrc4 0111
a8 vinrc4 a6 0111
a9 z55 z57 0110
a10 z53 a7 0111
a11 z53 z57 0110
a12 z51 a6 0001
a14 z53 a9 0100
a15 vinrc4 a9 0010
a16 z51 a14 0100
a17 vinrc4 a14 0010
a18 z51 z53 0110
a19 vinrc4 a12 0111
a20 a11 a15 0100
a21 a11 a18 0010
a22 a9 a18 0001
a23 a17 a22 0010
a24 a18 a20 0100
a25 vinrc4 a16 0010
a26 a19 a22 0111
a27 a15 a21 0010
a28 z51 a10 0111
a29 a7 a21 0111
vinrc4 z56 z50 0111
vinrc5 z57 vinrc4 0100
vinrc5 a24 a20 a27 a15 a23 a17 a25 vinrc4 a19 a8 a26 a7 a29 a10 a28