3 2 1
x1 x2 x3 
z0 x1 x2 0001
z1 z0 x3 0001
z1 