8 35 8
x1 x2 x3 x4 x5 x6 x7 x8
z0 x1 x2 0110
z1 x2 x3 0110
z2 z0 z1 0111
z3 z0 x3 0110
z4 z2 z3 0110
z5 x4 z3 0110
z6 x4 x5 0110
z7 z5 z6 0010
z8 z3 z6 0110
z9 z2 z7 0110
z10 z4 z9 0010
z11 z8 x6 0110
z12 z11 x7 0110
z13 z8 x6 0001
z14 z11 x7 0001
z15 z13 z14 0110
z16 z12 x8 0110
z17 z12 x8 0001
z18 z9 z15 0110
z19 z18 z17 0110
z20 z9 z15 0001
z21 z18 z17 0001
z22 z20 z21 0110
z23 z10 z22 0110
a5 z19 z23 0110
a6 pufaj4 a5 0111
a7 z16 z23 0110
a8 a5 a7 0001
a9 a6 a7 0111
a11 pufaj4 a5 0010
a12 pufaj4 a8 0010
a13 a8 a12 0110
a14 a7 a11 0100
pufaj4 z23 z10 0111
pufaj5 z22 z10 0001
pufaj5 a14 a11 a12 pufaj4 a13 a6 a9