6 12 1
x1 x2 x3 x4 x5 x6 
z0 x1 x2 0110
z1 x3 x4 0110
z2 x1 x5 0110
z3 x3 x5 0110
z4 x2 x6 0110
z5 z1 z2 0110
z6 z1 z3 0111
z7 z0 z6 0110
z8 z5 z6 0100
z9 z4 z7 0100
z10 z4 z8 0110
z11 z9 z10 1000
z11 