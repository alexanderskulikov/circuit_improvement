6 11 1
x1 x2 x3 x4 x5 x6
a3 x2 x3 1001
a4 x3 x1 1001
a5 x1 a3 1001
a6 a3 a4 1110
c3 x5 x6 1001
c4 x6 x4 1001
c5 x4 c3 1001
c6 c3 c4 1110
d1 a5 c5 0110
d2 a6 c6 1001
d3 d1 d2 0001
d3