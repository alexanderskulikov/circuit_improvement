4 6 1
x1 x2 x3 x4
b5 x3 x1 1000
c5 x2 x1 0100
d5 x2 x3 1101
d6 x4 d5 1011
d7 c5 d6 0100
d8 b5 d7 1001
d8