10 31 4
x0 x1 x2 x3 x4 x5 x6 x7 x8 x9
z0 x2 x3 0110
z1 x4 x5 0110
z2 x6 x7 0110
z3 x8 x9 0110
z4 x0 x1 0110
z5 x0 x1 0001
z6 x2 z4 0110
z7 z0 z6 0111
z8 z0 z4 0110
z9 z7 z8 0110
z10 x4 z8 0110
z11 z8 z1 0110
z12 z10 z1 0010
z13 z7 z12 0110
z14 x6 z11 0110
z15 z2 z14 0111
z16 z2 z11 0110
z17 z15 z16 0110
z18 x8 z16 0110
z19 z16 z3 0110
z20 z18 z3 0010
z21 z15 z20 0110
z22 z9 z5 0110
z23 z13 z22 0111
z24 z13 z5 0110
z25 z23 z24 0110
z26 z17 z24 0110
z27 z24 z21 0110
z28 z26 z21 0010
z29 z23 z28 0110
z30 z25 z29 0010
z19 z27 z29 z30