6 23 6
x1 x2 x3 x4 x5 x6
z0 x1 x2 0110
z1 x2 x3 0110
z2 z0 z1 0111
z3 z0 x3 0110
z4 z2 z3 0110
z5 x4 z3 0110
z6 x4 x5 0110
z7 z5 z6 0010
z8 z3 z6 0110
z9 z2 z7 0110
z11 z8 x6 0110
z12 z8 x6 0001
z13 z9 z12 0110
z14 z9 z12 0001
a3 z11 pntcy5 0111
a4 z11 pntcy5 0001
a5 z13 pntcy5 0001
a6 a4 a5 0110
a8 z13 pntcy5 0111
a9 a3 a8 0001
a10 z11 a8 0111
pntcy4 z4 z9 0010
pntcy5 z14 pntcy4 0110
a5 a6 pntcy5 a9 a8 a10