10 45 10
x1 x2 x3 x4 x5 x6 x7 x8 x9 x10
z0 x2 x3 0110
z1 x1 x2 0110
z2 x3 z1 0110
z3 x4 z2 0110
z4 x4 x5 0110
z5 z3 z4 0010
z6 z4 z2 0110
z7 z0 z1 0111
z8 z5 z7 0110
z9 z6 x6 0110
z10 z6 x6 0001
z11 z8 z10 0110
z12 z8 z10 0001
z13 z9 x7 0110
z14 x7 x8 0110
z15 z13 z14 0111
z16 z13 x8 0110
z17 z15 z16 0110
z18 x9 z16 0110
z19 x9 x10 0110
z20 z18 z19 0010
z21 z16 z19 0110
z22 z15 z20 0110
z23 z17 z22 0010
z24 z22 z11 0110
z25 z22 z11 0001
z26 z23 z25 0110
z27 z26 z12 0110
z28 z7 z2 0110
z29 z8 z28 1011
z30 z27 z29 1001
a6 z21 z24 0110
a7 cllyy5 a6 0010
a8 z30 a6 0001
a10 cllyy3 cllyy5 0001
a11 cllyy3 a7 0111
a12 a8 a10 0100
a13 a6 a11 0111
a14 a8 a10 0111
a15 cllyy5 a11 0111
a16 z24 cllyy4 0001
a17 a7 a12 0100
cllyy3 z26 z30 0111
cllyy4 z30 cllyy3 0100
cllyy5 z24 cllyy4 0111
a16 a17 cllyy4 a12 a10 a14 cllyy3 a11 a15 a13