4 3 1
a b c d
e1 b d 0001
e2 a e1 0111
e3 e2 c 0111
e3