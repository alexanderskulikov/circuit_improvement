2 1 1
x1 x2
z1 x1 x2 0001
z1 