5 8 1
z12 z16 z18 x8 x9
5 z18 x8 0110
6 z12 z16 0110
7 z16 x9 0110
8 z16 z18 0110
9 5 6 0010
10 7 8 0100
11 9 10 0001
12 z18 11 0110
12