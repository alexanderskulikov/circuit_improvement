6 13 1
x1 x2 x3 x4 x5 x6
z1 x2 x3 0110
c5 x2 x1 0110
c6 z1 c5 0111
d5 x3 c5 0110
z5 x4 d5 0110
z6 x4 x5 0110
z7 z5 z6 0010
c7 z7 c6 0110
e5 c7 z6 1101
e6 c6 e5 1110
e7 d5 e6 0110
e8 x6 c7 1110
e9 e7 e8 1110
e9