5 11 1
x1 x2 x3 x4 x5 
z0 x1 x2 1001
z1 x3 x4 0110
z2 x3 x4 0001
z3 x2 z1 0001
z4 z0 z1 1001
z5 z2 z3 0110
z6 x1 z5 0110
z7 z4 z6 1011
z8 x5 z7 1000
z9 z7 z5 1101
z10 z8 z9 0110
z10 