4 6 1
a b c d
m10 c b 1110
n5 m10 d 1011
n6 b d 0111
n7 a n5 0100
n8 c n6 0111
n9 n7 n8 0100
n9