3 5 2
x1 x2 x3
b3 x2 x3 0111
b4 x2 x3 1110
b5 x1 b3 1110
b6 x1 b3 0111
b7 b4 b5 1110
b7 b6