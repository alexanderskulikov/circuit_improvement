4 9 1
x1 x2 x3 x4
t1 x1 x2 0110
t2 x1 x2 1110
z0 t1 t2 0110
z1 t1 t2 0001
z2 z1 x4 1001
z3 x3 z0 0110
z4 z2 x3 1001
z5 z1 z3 0100
z6 z4 z5 1000
z6