4 5 1
a b c d
f4 b c 1001
f5 d f4 1001
f6 b f4 1011
f7 a f6 1110
f8 f5 f7 1011
f8