11 31 1
x1 x2 x3 x4 x5 x6 x7 x8 x9 x10 x11
z0 x1 x2 0110
z3 z0 x3 0001
z5 x4 x5 0110
z6 x6 x7 0110
z7 x4 s6 0110
s6 x3 z0 0110
z10 y5 s7 0110
s7 z5 s6 0110
z11 x6 s7 0110
z13 z11 z6 0010
z15 x8 x9 0110
z16 x10 x11 0110
z17 x8 s8 0110
s8 z6 s7 0110
z18 z15 z17 0111
z20 z18 s9 0110
s9 z15 s8 0110
z21 x10 s9 0110
z23 z21 z16 0010
z24 z18 z23 0110
z27 y6 j7 0110
j7 z3 j6 0111
j6 x2 x1 0001
z29 z20 z27 0110
q7 z27 y8 0110
j8 z10 j7 0110
p5 z24 z29 0111
y5 z7 z5 0111
y6 z13 y5 0110
y7 j8 y6 0111
y8 p5 y7 0001
q7