3 4 1
x1 x2 x3 
z0 x1 x2 0001
z1 x1 x2 1000
z2 x3 z1 0010
z3 z0 z2 0111
z3 