10 34 4
x1 x2 x3 x4 x5 x6 x7 x8 x9 x10 
z0 x1 x2 0110
z1 x2 x3 0110
z2 z0 z1 0111
z3 z0 x3 0110
z4 z2 z3 0110
z5 x4 z3 0110
z6 x4 x5 0110
z7 z5 z6 0010
z8 z3 z6 0110
z9 z2 z7 0110
z10 z4 z9 0010
z11 z8 x6 0110
z12 z8 x6 0001
z13 z9 z12 0110
z14 z9 z12 0001
z15 z10 z14 0110
z16 z11 x7 0110
z17 x7 x8 0110
z18 z16 z17 0111
z19 z16 x8 0110
z20 z18 z19 0110
z21 x9 z19 0110
z22 x9 x10 0110
z23 z21 z22 0010
z24 z19 z22 0110
z25 z18 z23 0110
z26 z20 z25 0010
z27 z25 z13 0110
z28 z25 z13 0001
z29 z15 z26 0110
z30 z26 z28 0110
z31 z29 z30 0111
z32 z29 z28 0110
z33 z31 z32 0110
z24 z27 z32 z33 