14 48 4
x1 x2 x3 x4 x5 x6 x7 x8 x9 x10 x11 x12 x13 x14
z0 x3 x4 0110
z1 x5 x6 0110
z2 x7 x8 0110
z3 x9 x10 0110
z4 x11 x12 0110
z5 x13 x14 0110
z6 x1 x2 0110
z7 x1 x2 0001
z8 x3 z6 0110
z9 z0 z8 0111
z10 z0 z6 0110
z11 z9 z10 0110
z12 x5 z10 0110
z13 z10 z1 0110
z14 z12 z1 0010
z15 z9 z14 0110
z16 x7 z13 0110
z17 z2 z16 0111
z18 z2 z13 0110
z19 z17 z18 0110
z20 x9 z18 0110
z21 z18 z3 0110
z22 z20 z3 0010
z23 z17 z22 0110
z24 x11 z21 0110
z25 z4 z24 0111
z26 z4 z21 0110
z27 z25 z26 0110
z28 x13 z26 0110
z29 z26 z5 0110
z30 z28 z5 0010
z31 z25 z30 0110
z32 z11 z7 0110
z33 z15 z32 0111
z34 z15 z7 0110
z35 z33 z34 0110
z36 z19 z34 0110
z37 z34 z23 0110
z38 z36 z23 0010
z39 z33 z38 0110
z40 z37 z31 0110
z41 z27 z31 0010
z42 z37 z31 0001
z43 z41 z42 0110
z44 z43 z39 0110
z45 z35 z39 0010
z46 z43 z39 0001
z47 z45 z46 0110
z29 z40 z44 z47