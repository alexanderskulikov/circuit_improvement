3 4 1
x1 x2 x3 
z1 x1 x2 0110
z2 x3 x2 0110
z3 z2 z1 0100
z4 x1 z3 0110
z4