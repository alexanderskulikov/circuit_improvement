12 31 1
x1 x2 x3 x4 x5 x6 x7 x8 x9 x10 x11 x12
z1 x1 x2 0001
z2 x1 x2 0111
z3 z2 x3 0001
z4 z2 x3 0111
z5 z4 x4 0001
z6 z4 x4 0111
z7 z6 x5 0001
z8 z6 x5 0111
z9 z8 x6 0001
z10 z8 x6 0111
z11 z10 x7 0001
z12 z10 x7 0111
z13 z12 x8 0001
z14 z12 x8 0111
z15 z14 x9 0001
z16 z14 x9 0111
z17 z16 x10 0001
z18 z16 x10 0111
z19 z18 x11 0001
z20 z18 x11 0111
z21 z20 x12 0001
z22 z1 z3 0111
z23 z22 z5 0111
z24 z23 z7 0111
z25 z24 z9 0111
z26 z25 z11 0111
z27 z26 z13 0111
z28 z27 z15 0111
z29 z28 z17 0111
z30 z29 z19 0111
z31 z30 z21 0111
z31