7 16 1
x1 x2 x3 x4 x5 x6 x7
z0 x1 x2 1001
z1 x1 x2 1000
z2 z1 x3 1001
z3 z0 z2 1001
z4 z1 z3 0100
z5 x4 z2 1001
z6 z5 z4 0111
z7 z6 x5 0110
z8 z7 z4 0110
z9 z8 x4 0110
z10 z9 z6 0001
z11 z10 x6 1001
z12 z7 z11 1001
z13 z10 z12 0100
z14 x7 z11 0110
z15 z13 z14 0100
z15