11 55 11
x1 x2 x3 x4 x5 x6 x7 x8 x9 x10 x11
z0 x1 x2 0110
z1 z0 x3 0110
z2 x1 x2 0001
z3 z0 x3 0001
z4 z2 z3 0110
z5 x4 x5 0110
z6 x6 x7 0110
z7 x4 z1 0110
z8 z5 z7 0111
z9 z5 z1 0110
z10 z8 z9 0110
z11 x6 z9 0110
z12 z9 z6 0110
tmpneg1 z6 z6 1100
z13 z11 tmpneg1 0001
z14 z8 z13 0110
z15 x8 x9 0110
z16 x10 x11 0110
z17 x8 z12 0110
z18 z15 z17 0111
z19 z15 z12 0110
z20 z18 z19 0110
z21 x10 z19 0110
z22 z19 z16 0110
tmpneg2 z16 z16 1100
z23 z21 tmpneg2 0001
z24 z18 z23 0110
z25 z10 z4 0110
z26 z14 z25 0111
z27 z14 z4 0110
z29 z20 z27 0110
z30 z27 z24 0110
tmpneg3 z24 z24 1100
z31 z29 tmpneg3 0001
z32 z26 z31 0110
a4 z32 blzee4 0110
a5 z22 z30 0001
a6 z22 z30 0110
a7 blzee4 a6 0001
a8 blzee4 a5 0001
a9 a7 a8 0110
a10 z30 a4 0001
a12 a4 a5 0111
a13 blzee4 a10 0111
a14 z32 a6 0001
tmpneg4 z32 z32 1100
a15 tmpneg4 a10 0001
tmpneg5 a14 a14 1100
a16 a13 tmpneg5 0001
a17 z30 a12 0111
a18 a14 a16 0111
a19 a6 a17 0111
blzee3 z27 z26 0110
tmpneg6 z32 z32 1100
blzee4 tmpneg6 blzee3 0001
a8 a15 a9 blzee4 a16 a13 a18 a4 a12 a17 a19