4 6 1
x1 x2 x3 x4 
z0 x1 x2 1011
z1 x3 z0 1011
z2 x1 z1 1001
z3 x4 z0 0110
z4 x3 z3 0110
z5 z4 z2 0010
z5 