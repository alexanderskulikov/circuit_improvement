7 19 3
x1 x2 x3 x4 x5 x6 x7 
z0 x1 x2 0110
z1 x2 x3 0110
z2 z0 z1 0111
z3 z0 x3 0110
z5 x4 z3 0110
z6 x4 x5 0110
z10 a9 a10 0010
z11 a8 x6 0110
z12 x6 x7 0110
z13 z11 z12 0111
z14 z11 x7 0110
z15 z13 z14 0110
z16 a10 z15 0110
z17 a10 z15 0001
a6 z6 z5 1011
a7 z17 z10 0111
a8 z6 z3 0110
a9 z3 z2 0110
a10 z2 a6 1001
z14 z16 a7