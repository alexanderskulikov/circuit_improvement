3 3 1
x1 x2 x3 
z0 x2 x1 1101
z1 x3 z0 0100
z2 x1 z1 0110
z2 