4 5 1
x1 x2 x3 x4 
z0 x1 x4 1001
z1 x3 x2 0110
z2 z0 x3 1001
z3 x1 z1 0100
z4 z2 z3 1000
z4 