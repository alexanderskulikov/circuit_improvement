5 9 2
x1 x2 x3 x4 x5 
z0 x3 x2 1001
z1 z0 x1 0111
z2 z1 x4 0110
z3 z2 x1 0110
z4 z3 x3 0110
z5 z4 z1 0001
z6 z5 x5 1001
z7 z2 z6 1001
z8 z5 z7 0100
z8 z6 