4 8 2
a b c d
h6 b c 0001
h7 e9 h6 0111
e4 b d 0001
e5 c e4 0111
e6 a e5 0001
e7 a e5 0111
e8 b d 1001
e9 e6 e8 1011
e7 h7