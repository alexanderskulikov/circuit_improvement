2 1 1
x1 x2 
z0 x1 x2 0111
z0 