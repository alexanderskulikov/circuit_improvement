4 7 1
x1 x2 x3 x4 
z0 x1 x2 0001
z1 x3 x4 0110
z2 z0 z1 0001
z3 x1 x2 0110
z4 x3 x4 0001
z5 z3 z4 0001
z6 z2 z5 0111
z6 