5 10 1
x1 x2 x3 x4 x5
a2 e5 x3 0001
a3 e6 x4 0001
a4 e7 x5 0001
c2 a3 a4 0111
d5 x2 x1 0001
d6 c2 d5 1000
d7 a2 d6 1011
e5 x2 x1 0111
e6 x3 e5 0111
e7 x4 e6 0111
d7