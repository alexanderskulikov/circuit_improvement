3 5 2
a b c
e1 b c 0110
e2 b c 0001
e3 e2 a 0001
e4 e1 e3 0111
e5 a e2 0111
e5 e4