4 7 1
x1 x2 x3 x4
z0 x1 x2 1001
z1 x1 x2 1000
z2 z1 x3 1001
z3 z0 z2 1001
z4 z1 z3 0100
z5 x4 z2 0110
z6 z4 z5 0100
z6