2 2 2
x1 x2 
z0 x1 x2 0110
z1 x1 x2 0001
z0 z1 