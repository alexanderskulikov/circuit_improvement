5 9 1
x1 x2 x3 x4 x5
z1 x1 x2 0110
z2 x2 x3 0110
z3 x3 z1 1001
z4 z2 z1 1000
z5 x4 z3 0110
z6 x4 x5 0110
z7 z5 z6 0010
z8 z7 z4 1000
z9 z8 z3 1001
z9