3 3 1
x1 x2 x3
z0 x2 x3 1001
z1 x1 x2 0110
z2 z0 z1 0010
z2