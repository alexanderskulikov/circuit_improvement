7 16 2
x1 x2 x3 x4 x5 x6 x7 
z0 x3 x2 1001
z1 z0 x1 0111
z2 z1 x4 0110
z3 z2 x1 0110
z4 z3 x3 0110
z5 z4 z1 0001
z6 z5 x5 1001
z7 z2 z6 1001
z8 z5 z7 0100
z9 z6 z8 0010
z10 x7 z9 1001
z11 x6 z10 0110
z12 x6 z9 1000
z13 z8 z12 0110
z14 x7 z13 1001
z15 z11 z13 0010
z15 z14 