7 17 1
x1 x2 x3 x4 x5 x6 x7 
z0 x1 x2 0110
z1 x2 x3 0110
z2 z0 z1 0111
z3 z0 x3 0110
z4 z2 z3 0110
z5 x4 z3 0110
z6 x4 x5 0110
z7 z5 z6 0010
z8 z3 z6 0110
z9 z2 z7 0110
z10 z4 z9 0010
z16 z9 a6 0001
z17 z10 z16 0110
a3 x7 z8 0001
a4 x7 z8 1000
a5 x6 a4 0010
a6 a3 a5 0111
z17 