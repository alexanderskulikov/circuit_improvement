7 19 3
x1 x2 x3 x4 x5 x6 x7
z0 x1 x2 0110
z1 x2 x3 0110
z3 z0 x3 0110
z5 z3 x4 0110
z6 x4 x5 0110
z8 z5 x5 0110
z10 z8 x6 0110
z11 x6 x7 0110
z12 z10 z11 0111
z13 z10 x7 0110
z14 z12 z13 0110
z16 7 z14 0110
z17 9 z16 0111
z18 9 z14 0110
z19 z17 z18 0110
6 z5 z6 0010
7 z3 6 0110
8 z0 z1 0111
9 6 8 0110
z13 z18 z19