6 12 1
x1 x2 x3 x4 x5 x6
z0 x2 x1 1001
z1 z0 x3 0110
z2 x2 z1 0110
z3 z2 z0 0001
z4 z3 x4 1001
z5 z1 z4 1001
z6 z3 z5 0100
z7 z6 x6 1001
z8 x5 z4 0110
z9 z7 x5 1001
z10 z6 z8 0100
z11 z9 z10 1000
z11