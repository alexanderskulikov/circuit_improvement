4 8 2
a b c d
g6 g4 g5 1101
g3 c b 1001
g4 c b 1110
g5 d g3 0010
h5 g6 a 1110
h6 d g3 0110
h7 g6 a 0111
h8 h5 h6 1110
h7 h8