5 10 1
x1 x2 x3 x4 x5
z0 x1 x2 1001
z1 x1 x2 1000
z2 z1 x3 1001
z3 z0 z2 1001
z4 z1 z3 0100
z5 z4 x5 1001
z6 x4 z2 0110
z7 z5 x4 1001
z8 z4 z6 0100
z9 z7 z8 1000
z9