13 46 1
x1 x2 x3 x4 x5 x6 x7 x8 x9 x10 x11 x12 x13
z0 x1 x2 0110
z1 x2 x3 0110
z2 z0 z1 0111
z3 z0 x3 0110
z4 z2 z3 0110
z5 x4 z3 0110
z6 x4 x5 0110
z7 z5 z6 0010
z8 z3 z6 0110
z9 z2 z7 0110
z10 z4 z9 0010
z11 z8 x6 0110
z12 z11 x7 0110
z13 z8 x6 0001
z14 z11 x7 0001
z15 z13 z14 0110
z16 z9 z15 0110
z17 z9 z15 0001
z18 z10 z17 0110
z19 z12 x8 0110
z20 x8 x9 0110
z21 z19 z20 0111
z22 z19 x9 0110
z23 z21 z22 0110
z24 x10 z22 0110
z25 x10 x11 0110
z26 z24 z25 0010
z27 z22 z25 0110
z28 z21 z26 0110
z29 z23 z28 0010
z30 z27 x12 0110
z31 z30 x13 0110
z32 z27 x12 0001
z33 z30 x13 0001
z34 z32 z33 0110
z35 z28 z34 0110
z36 z28 z34 0001
z37 z29 z36 0110
z38 z16 z35 0110
z39 z16 z35 0001
z40 z18 z37 0110
z42 z18 z37 0001
z45 z31 z38 0001
t4 z45 z39 0110
t5 z40 t4 0001
t6 z42 t5 0111
t6