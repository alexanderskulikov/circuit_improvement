10 32 4
x1 x2 x3 x4 x5 x6 x7 x8 x9 x10 
z0 x2 x3 0110
z1 x1 x2 0110
z2 x3 z1 0110
z3 x4 z2 0110
z4 x4 x5 0110
z5 z3 z4 0010
z6 z4 z2 0110
z7 z0 z1 0111
z8 z5 z7 0110
z9 z6 x6 0110
z10 z6 x6 0001
z11 z8 z10 0110
z12 z8 z10 0001
z13 z9 x7 0110
z14 x7 x8 0110
z15 z13 z14 0111
z16 z13 x8 0110
z17 z15 z16 0110
z18 x9 z16 0110
z19 x9 x10 0110
z20 z18 z19 0010
z21 z16 z19 0110
z22 z15 z20 0110
z23 z17 z22 0010
z24 z22 z11 0110
z25 z22 z11 0001
z26 z23 z25 0110
z27 z26 z12 0110
z28 z7 z2 0110
z29 z8 z28 1011
z30 z27 z29 1001
z31 z26 z30 0010
z21 z24 z30 z31 