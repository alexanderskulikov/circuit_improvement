4 7 1
x1 x2 x3 x4
z1 x1 x2 0110
z2 x2 x3 0110
z3 x3 z1 1001
z4 z2 z1 1000
z5 x4 z3 0100
z6 z4 z5 1000
z7 z6 z3 1001
z7