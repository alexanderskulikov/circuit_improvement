12 29 1
x1 x2 x3 x4 x5 x6 x7 x8 x9 x10 x11 x12
z0 x1 x2 0111
z1 z0 x3 0111
z2 z1 x4 0111
z3 x5 x6 0111
z4 z3 x7 0111
z5 z4 x8 0111
z6 x9 x10 0111
z7 z6 x11 0111
z8 z7 x12 0111
z9 x1 x5 0111
z10 z9 x9 0111
z11 x2 x6 0111
z12 z11 x10 0111
z13 x3 x7 0111
z14 z13 x11 0111
z15 x4 x8 0111
z16 z15 x12 0111
z17 z2 z5 0001
z18 z2 z5 0111
z19 z18 z8 0001
z20 z17 z19 0111
z21 z10 z12 0001
z22 z10 z12 0111
z23 z22 z14 0001
z24 z22 z14 0111
z25 z24 z16 0001
z26 z21 z23 0111
z27 z25 z26 0111
z28 z20 z27 0111
z28