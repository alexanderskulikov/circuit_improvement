14 68 14
x1 x2 x3 x4 x5 x6 x7 x8 x9 x10 x11 x12 x13 x14
z0 x3 x4 0110
z1 x5 x6 0110
z2 x7 x8 0110
z3 x9 x10 0110
z4 x11 x12 0110
z5 x13 x14 0110
z6 x1 x2 0110
z7 x1 x2 0001
z8 x3 z6 0110
z9 z0 z8 0111
z10 z0 z6 0110
z11 z9 z10 0110
z12 x5 z10 0110
z13 z10 z1 0110
z14 z12 z1 0010
z15 z9 z14 0110
z16 x7 z13 0110
z17 z2 z16 0111
z18 z2 z13 0110
z19 z17 z18 0110
z20 x9 z18 0110
z21 z18 z3 0110
z22 z20 z3 0010
z23 z17 z22 0110
z24 x11 z21 0110
z25 z4 z24 0111
z26 z4 z21 0110
z27 z25 z26 0110
z28 x13 z26 0110
z29 z26 z5 0110
z30 z28 z5 0010
z31 z25 z30 0110
z32 z11 z7 0110
z33 z15 z32 0111
z34 z15 z7 0110
z35 z33 z34 0110
z36 z19 z34 0110
z37 z34 z23 0110
z38 z36 z23 0010
z39 z33 z38 0110
z40 z37 z31 0110
z41 z27 z31 0010
z42 z37 z31 0001
z43 z41 z42 0110
z44 z43 z39 0110
z46 z43 z39 0001
a4 z40 ghujg5 0001
a5 z44 ghujg5 0111
a6 z44 a4 0001
a7 z40 z44 0001
a8 z29 a4 0110
a9 z40 a5 0111
a10 z44 ghujg5 0001
a11 z29 a7 0001
a13 a11 ghujg5 0111
a14 z29 a9 0111
a15 a7 a13 0111
a16 z29 a5 0111
a17 a8 a10 0001
a18 a9 a16 0001
a19 a5 a8 0001
a20 a15 a19 0111
a21 a4 a10 0111
a22 z44 a19 0100
a23 a21 a22 0010
a24 a21 a22 0111
ghujg4 z39 z35 0100
ghujg5 z46 ghujg4 0110
a6 a17 a10 a23 a21 a24 ghujg5 a13 a15 a20 a5 a18 a9 a14