5 9 1
x1 x2 x3 x4 x5
g4 x4 x3 1011
j8 k6 x3 1001
k6 x4 x2 1001
m6 x5 x1 0010
m7 k6 m6 0110
m8 x5 g4 0001
m9 x1 m8 0010
m10 j8 m9 0110
m11 m7 m10 0001
m11