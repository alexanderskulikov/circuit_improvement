5 10 1
x1 x2 x3 x4 x5
z0 x1 x2 0110
z1 x1 x2 0001
z2 x3 z0 1001
z3 z2 z1 0111
z4 x4 z3 0110
z5 z4 z1 0110
z6 z5 x3 0110
z7 z6 z3 0001
z8 x5 z4 1001
z9 z7 z8 1000
z9