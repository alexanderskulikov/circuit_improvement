5 12 3
x1 x2 x3 x4 x5 
z0 x1 x2 0110
z1 x2 x3 0110
z2 z0 z1 0111
z3 z0 x3 0110
z4 z2 z3 0110
z5 z3 x4 0110
z6 x4 x5 0110
z7 z5 z6 0111
z8 z5 x5 0110
z9 z7 z8 0110
z10 z4 z9 0110
z11 z4 z9 0001
z8 z10 z11 