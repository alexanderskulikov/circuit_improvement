4 7 1
x1 x2 x3 x4 
z4 x1 x2 0111
a5 x1 x2 0110
a6 x4 z4 1001
a7 x3 a6 0010
a8 x4 a5 0111
a9 a6 a8 0110
a10 a7 a9 1011
a10