3 3 1
x1 x2 x3 
z0 x3 x1 1001
z1 x2 x1 0111
z2 z0 z1 0100
z2 