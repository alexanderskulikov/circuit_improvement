3 4 1
x1 x2 x3
z0 x1 x2 0110
z1 x1 x2 0001
z2 x3 z0 0110
z3 z1 z2 0100
z3