11 34 4
x1 x2 x3 x4 x5 x6 x7 x8 x9 x10 x11
z0 x1 x2 0110
z1 z0 x3 0110
z2 x1 x2 0001
z3 z0 x3 0001
z4 z2 z3 0110
z5 x4 x5 0110
z6 x6 x7 0110
z7 x4 z1 0110
z8 z5 z7 0111
z9 z5 z1 0110
z10 z8 z9 0110
z11 x6 z9 0110
z12 z9 z6 0110
z13 z11 z6 0010
z14 z8 z13 0110
z15 x8 x9 0110
z16 x10 x11 0110
z17 x8 z12 0110
z18 z15 z17 0111
z19 z15 z12 0110
z20 z18 z19 0110
z21 x10 z19 0110
z22 z19 z16 0110
z23 z21 z16 0010
z24 z18 z23 0110
z25 z10 z4 0110
z26 z14 z25 0111
z27 z14 z4 0110
z28 z26 z27 0110
z29 z20 z27 0110
z30 z27 z24 0110
z31 z29 z24 0010
z32 z26 z31 0110
z33 z28 z32 0010
z22 z30 z32 z33