6 13 3
x1 x2 x3 x4 x5 x6
z0 x1 x2 0110
z2 a5 x4 0110
a5 x3 z0 0110
z4 b10 x6 0110
z10 x1 z0 0010
a6 z10 a5 0110
a7 z2 a6 0111
b6 x5 a5 1101
b7 z4 b6 1011
b8 a7 b7 1000
b9 x5 b8 0001
b10 z2 x5 0110
b11 x3 b8 1011
z4 b11 b9