7 18 1
x1 x2 x3 x4 x5 x6 x7
z0 x1 x2 0110
z1 x2 x3 0110
z3 z0 x3 0110
z4 b5 z3 0110
b5 z0 z1 0111
z5 x4 z3 0110
z6 x4 x5 0110
z8 z3 z6 0110
z10 z4 c7 0010
z11 z8 x6 0110
z12 x6 x7 0110
z13 z11 z12 0111
a7 z10 c9 1000
a8 c7 a7 1001
c6 z6 z5 0100
c7 b5 c6 0110
c8 x7 c7 0110
c9 z13 c8 0100
a8