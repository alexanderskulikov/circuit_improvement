7 17 1
x1 x2 x3 x4 x5 x6 x7
z0 x1 x2 0110
z1 x2 x3 0110
z2 z0 z1 0111
z3 z0 x3 0110
z5 z3 x4 0110
z6 x4 x5 0110
z8 z5 x5 0110
z10 z8 x6 0110
b5 x7 z10 0110
a7 z3 a5 1001
a5 z6 z5 1011
a6 z2 a5 1001
c5 a7 a6 0010
d6 c5 e7 0100
e5 z10 x6 1011
e6 a6 e5 1001
e7 b5 e6 0001
d6