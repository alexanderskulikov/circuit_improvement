5 12 1
xx1 xx2 x3 x4 x5
x1 xx1 xx2 0110
x2 xx1 xx2 1110
s5 x1 x2 0110
s6 x3 s5 0110
s7 x1 x4 0110
s8 x4 x5 0110
s9 x2 x3 0001
s10 s7 s9 0110
s11 s6 s9 1101
s12 s8 s11 0110
s13 s8 s10 1000
s14 s12 s13 0010
s14 