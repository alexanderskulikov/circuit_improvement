5 13 2
a b c d x
g6 g4 g5 1101
g3 c b 1001
g4 c b 1110
g5 d g3 0010
h5 g6 a 1110
h6 d g3 0110
h7 g6 a 0111
h8 h5 h6 1110
e1 h8 x 0110
e2 h8 x 0001
e3 e2 h7 0001
e4 e1 e3 0111
e5 h7 e2 0111
e5 e4