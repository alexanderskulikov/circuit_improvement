4 7 2
x1 x2 x3 x4 
z0 x2 x1 0010
z1 x4 z0 1001
z2 x3 z1 0110
z3 x3 z0 1000
z4 x1 z3 0110
z5 x4 z4 1001
z6 z2 z4 0010
z6 z5 