5 8 1
x1 x2 x3 x4 x5 
z0 x3 x2 1001
z1 z0 x1 0111
z2 x4 z1 0110
z3 z2 x1 0110
z4 z3 x3 0110
z5 z4 z1 0001
z6 x5 z2 1001
z7 z5 z6 1000
z7 