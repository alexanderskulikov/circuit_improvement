5 9 1
x1 x2 x3 x4 x5
z1 x2 x3 0110
z3 b5 x3 0110
b5 x1 x2 0110
z5 z3 x4 0110
z8 z5 x5 0110
e5 z1 b5 0111
e6 x4 z5 1110
e7 e5 e6 1001
d7 z8 e7 0100
d7