4 6 1
x1 x2 x3 x4
z0 x1 x2 0110
z1 x3 x4 0110
z2 x1 x3 0110
z3 z1 z2 0111
z4 z0 z3 0100
z5 z1 z4 0110
z5