3 4 2
x1 x2 x3 
z0 x2 x1 1000
z1 x3 z0 0010
z2 x3 z0 1001
z3 x1 z1 0110
z3 z2 