4 7 1
x1 x2 x3 x4 
z0 x1 x2 0001
z1 x3 x4 0111
z2 x3 x4 0001
z3 x1 z2 1000
z4 x2 z3 1011
z5 z1 z4 1110
z6 z0 z5 1011
z6 