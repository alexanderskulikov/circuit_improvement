3 4 1
x1 x2 x3
z3 x1 x3 1000
z4 x2 z3 0111
z5 x3 z4 0110
z6 x1 z5 1001
z6