13 43 4
x1 x2 x3 x4 x5 x6 x7 x8 x9 x10 x11 x12 x13
z0 x6 x7 0110
z1 x8 x9 0110
z2 x10 x11 0110
z3 x12 x13 0110
z4 x1 x2 0110
z5 x2 x3 0110
z6 z4 z5 0111
z7 z4 x3 0110
z8 z6 z7 0110
z9 x4 z7 0110
z10 x4 x5 0110
z11 z9 z10 0010
z12 z7 z10 0110
z13 z6 z11 0110
z14 z8 z13 0010
z15 x6 z12 0110
z16 z0 z15 0111
z17 z0 z12 0110
z18 z16 z17 0110
z19 x8 z17 0110
z20 z17 z1 0110
z21 z19 z1 0010
z22 z16 z21 0110
z23 x10 z20 0110
z24 z2 z23 0111
z25 z2 z20 0110
z26 z24 z25 0110
z27 x12 z25 0110
z28 z25 z3 0110
z29 z27 z3 0010
z30 z24 z29 0110
z31 z18 z13 0110
z32 z22 z31 0111
z33 z22 z13 0110
z34 z32 z33 0110
z35 z26 z33 0110
z36 z33 z30 0110
z37 z35 z30 0010
z38 z32 z37 0110
z39 z14 z38 0110
z40 z34 z38 0010
z41 z14 z38 0001
z42 z40 z41 0110
z28 z36 z39 z42