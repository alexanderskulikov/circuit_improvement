7 18 1
x1 x2 x3 x4 x5 x6 x7
z0 x1 x2 0110
z1 x2 x3 0110
z3 z0 x3 0110
z5 z3 x4 0110
z6 x4 x5 0110
z8 z5 x5 0110
z11 x6 x7 0110
c5 x6 z8 0110
a7 z3 a6 1001
a6 z6 z5 1011
a8 z1 z0 0111
b6 d5 a7 0100
b9 b6 d8 1011
c6 z11 c5 1000
d5 a6 a8 1001
d6 c6 x7 0010
d7 c6 d5 1000
d8 d6 d7 0111
b9