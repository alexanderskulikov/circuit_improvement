6 15 3
x1 x2 x3 x4 x5 x6 
z0 x1 x2 0110
z1 x3 z0 0110
z2 x4 z1 0110
z3 x5 z2 0110
z4 x6 z3 0110
z5 x1 x2 0001
z6 x3 z5 0001
z7 x4 z6 0001
z8 x5 z7 0001
z9 x6 z8 0001
z10 x1 x2 0111
z11 x3 z10 0111
z12 x4 z11 0111
z13 x5 z12 0111
z14 x6 z13 0111
z4 z9 z14 