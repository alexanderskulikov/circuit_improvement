10 44 10
x0 x1 x2 x3 x4 x5 x6 x7 x8 x9
z0 x2 x3 0110
z1 x4 x5 0110
z2 x6 x7 0110
z3 x8 x9 0110
z4 x0 x1 0110
z5 x0 x1 0001
z6 x2 z4 0110
z7 z0 z6 0111
z8 z0 z4 0110
z9 z7 z8 0110
z10 x4 z8 0110
z11 z8 z1 0110
z12 z10 z1 0010
z13 z7 z12 0110
z14 x6 z11 0110
z15 z2 z14 0111
z16 z2 z11 0110
z17 z15 z16 0110
z18 x8 z16 0110
z19 z16 z3 0110
z20 z18 z3 0010
z21 z15 z20 0110
z22 z9 z5 0110
z23 z13 z22 0111
z24 z13 z5 0110
z26 z17 z24 0110
z27 z24 z21 0110
z28 z26 z21 0010
z29 z23 z28 0110
a4 z27 z29 0001
a7 z19 z27 0110
a8 z29 a7 0001
a9 arfvx6 a8 0111
a10 z19 z27 0001
a11 arfvx5 a7 0001
a12 z27 arfvx5 0001
a13 z29 arfvx6 0111
a14 a10 a13 0111
a15 a7 a14 0111
a16 z27 a14 0111
a17 arfvx6 a8 0010
arfvx4 z24 z23 0110
arfvx5 z29 arfvx4 0100
arfvx6 a4 arfvx5 0110
a12 a11 arfvx5 a17 arfvx6 a9 a13 a14 a16 a15