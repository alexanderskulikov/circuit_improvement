6 12 1
x1 x2 x3 x4 x5 x6 
z0 x3 x2 1001
z1 z0 x1 0111
z2 z1 x4 0110
z3 z2 x1 0110
z4 z3 x3 0110
z5 z4 z1 0001
z6 x5 z5 1001
z7 z2 z6 1001
z8 z5 z7 0100
z9 z8 z6 1000
z10 x6 z9 0010
z11 z8 z10 0110
z11 