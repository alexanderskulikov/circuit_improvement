5 9 1
x1 x2 x3 x4 x5
z5 x1 x2 0110
z6 x3 z5 0110
z7 x4 x5 0110
z8 x4 z6 0110
z9 x2 x3 0110
z10 z7 z8 0111
z11 z5 z9 0111
z12 z10 z11 0001
z13 z6 z12 0110
z13