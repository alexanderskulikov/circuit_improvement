5 14 2
x1 x2 x3 x4 x5
z0 x1 x2 0110
z1 x2 x3 0110
z2 z0 z1 0111
z3 z0 x3 0110
z4 z2 z3 0110
z5 z3 x4 0110
z6 x4 x5 0110
z7 z5 z6 0111
z8 z5 x5 0110
b3 z4 z7 0110
b4 z8 b3 0110
b5 z4 b4 0010
a1 b5 b4 0111
a3 b3 b5 0010
a1 a3