5 9 1
x1 x2 x3 x4 x5
a5 x1 a3 1001
z6 x4 x5 0110
a6 a3 a4 1110
a3 x2 x3 1001
a4 x3 x1 1001
b4 x4 z6 1000
b5 a6 b4 0110
b6 a5 z6 0110
b7 b5 b6 0001
b7