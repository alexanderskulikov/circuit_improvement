15 53 4
x1 x2 x3 x4 x5 x6 x7 x8 x9 x10 x11 x12 x13 x14 x15 
z0 x1 x2 0110
z1 x2 x3 0110
z2 z0 z1 0111
z3 z0 x3 0110
z4 z2 z3 0110
z5 x4 z3 0110
z6 x4 x5 0110
z7 z5 z6 0010
z8 z3 z6 0110
z9 z2 z7 0110
z10 z4 z9 0010
z11 z8 x6 0110
z12 x6 x7 0110
z13 z11 z12 0111
z14 z11 x7 0110
z15 z13 z14 0110
z16 z9 z15 0110
z17 z9 z15 0001
z18 z10 z17 0110
z19 z14 x8 0110
z20 x8 x9 0110
z21 z19 z20 0111
z22 z19 x9 0110
z23 z21 z22 0110
z24 x10 z22 0110
z25 x10 x11 0110
z26 z24 z25 0010
z27 z22 z25 0110
z28 z21 z26 0110
z29 z23 z28 0010
z30 z27 x12 0110
z31 x12 x13 0110
z32 z30 z31 0111
z33 z30 x13 0110
z34 z32 z33 0110
z35 z28 z34 0110
z36 z28 z34 0001
z37 z29 z36 0110
z38 z33 x14 0110
z39 x14 x15 0110
z40 z38 z39 0111
z41 z38 x15 0110
z42 z40 z41 0110
z43 z16 z35 0110
z44 z35 z42 0110
z45 z43 z44 0111
z46 z43 z42 0110
z47 z45 z46 0110
z48 z18 z37 0110
z49 z37 z47 0110
z50 z48 z49 0111
z51 z48 z47 0110
z52 z50 z51 0110
z41 z46 z51 z52 