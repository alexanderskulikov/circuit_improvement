6 22 6
a1 a2 a3 b1 b2 b3
x1 a1 b1 0001
x2 a2 b1 0001
x3 a3 b1 0001

y2 a1 b2 0001
y3 a2 b2 0001
y4 a3 b2 0001

z3 a1 b3 0001
z4 a2 b3 0001
z5 a3 b3 0001

-r2x x2 y2 0110
r3 x2 y2 0001

c1 x3 y3 0110
-c1 c1 r3 0110