4 6 1
x1 x2 x3 x4
f9 g8 g7 0100
g4 x2 x4 0110
g5 x4 x3 1001
g6 x2 x1 1001
g7 g5 g6 1001
g8 g4 g5 0100
f9