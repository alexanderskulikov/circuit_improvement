7 16 1
x1 x2 x3 x4 x5 x6 x7
z0 x1 x2 0110
z1 x1 x2 0001
z2 x3 z0 1001
z3 z2 z1 0111
z4 z3 x4 0110
z5 z4 z1 0110
z6 z5 x3 0110
z7 z6 z3 0001
z8 z7 x5 1001
z9 z4 z8 1001
z10 z7 z9 0100
z11 z10 x7 1001
z12 x6 z8 0110
z13 z11 x6 1001
z14 z10 z12 0100
z15 z13 z14 1000
z15