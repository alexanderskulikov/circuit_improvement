3 5 1
x1 x2 x3
t1 x1 x2 0110
t2 x1 x2 1110
z0 t2 x3 1001
z1 t1 t2 0110
z2 z0 z1 0010
z2