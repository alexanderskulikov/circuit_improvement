8 22 1
x1 x2 x3 x4 x5 x6 x7 x8
z0 x1 x2 0110
z1 x2 x3 0110
z2 z0 z1 0111
z3 z0 x3 0110
z5 x4 z3 0110
z6 x4 x5 0110
z7 z5 z6 0010
z8 z3 z6 0110
z9 z2 z7 0110
z12 z8 x6 0001
z13 z9 z12 0110
z14 z9 z12 0001
z17 x7 x8 0110
z22 b8 z13 0001
a5 z2 z3 0110
a6 z9 a5 0100
a7 z14 z22 0111
a8 a6 a7 0111
b5 z17 x7 1011
b6 z8 x6 1001
b7 z17 b6 1101
b8 b5 b7 0110
a8