6 13 1
x1 x2 x3 x4 x5 x6 
z0 x1 x2 0110
z1 x3 x4 0110
z2 x2 x5 0110
z3 z0 z2 1000
z4 x5 z3 0010
z5 z0 z4 0110
z6 x6 z5 0010
z7 z3 z6 0110
z8 z1 z7 0110
z9 x6 z5 0110
z10 x4 z9 0110
z11 z1 z10 1000
z12 z8 z11 1000
z12 