3 2 1
x1 x2 x3 
a3 x1 x2 0001
a4 a3 x3 0001
a4