6 15 1
x1 x2 x3 x4 x5 x6 
z0 x1 x2 1000
z1 x2 x3 0110
z2 x4 x5 1001
z3 x5 x6 1110
z4 x1 z1 1001
z5 x6 z2 1001
z6 x3 z4 1000
z7 z5 x4 0100
z8 z3 z7 1101
z9 z0 z8 0110
z10 z5 z9 1000
z11 z4 z10 1110
z12 z6 z0 0110
z13 z8 z12 0100
z14 z11 z13 0110
z14 