7 15 1
x1 x2 x3 x4 x5 x6 x7
z0 x2 x1 1001
z1 z0 x3 0110
z2 x2 z1 0110
z3 z2 z0 0001
z4 z3 x4 1001
z5 z1 z4 1001
z6 z3 z5 0100
z7 x5 z4 1001
z8 z7 z6 0111
z9 x6 z8 0110
z10 z9 z6 0110
z11 z10 x5 0110
z12 z11 z8 0001
z13 x7 z9 1001
z14 z12 z13 1000
z14