5 12 3
x1 x2 x3 x4 x5 
z0 x4 x2 1001
z1 x5 x1 1001
z2 x1 z0 0110
z3 z0 z1 1110
z4 x3 z2 0110
z5 z1 z4 0111
z6 x4 z3 0110
z7 z4 z6 1011
z8 x4 z7 1001
z9 z2 z8 1001
z10 x3 z1 1001
z11 z3 z5 1001
z9 z10 z11 