4 9 3
x1 x2 x3 x4 
z0 x1 x2 0110
z1 x2 x3 0110
z2 z0 z1 0111
z3 z0 x3 0110
z4 z2 z3 0110
z5 z3 x4 0110
z6 z3 x4 0001
z7 z4 z6 0110
z8 z4 z6 0001
z5 z7 z8 