3 5 2
x1 x2 x3 
z0 x1 x2 0110
z1 x2 x3 0110
z2 z0 z1 0111
z3 z0 x3 0110
z4 z2 z3 0110
z3 z4 