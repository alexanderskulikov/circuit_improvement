3 2 1
x1 x2 x3 
z0 x3 x2 0110
z1 x1 z0 0100
z1 