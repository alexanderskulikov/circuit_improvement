7 19 3
x1 x2 x3 x4 x5 x6 x7 
1899 1961 2001 0110
1961 x6 2000 0110
1937 1857 1998 1011
1857 x1 x3 0110
1896 x6 x7 0110
1957 x7 1919 0110
1919 x5 x4 1001
1941 2002 1978 1110
1978 1937 1976 1001
1959 x4 1999 1001
1976 1919 1959 0010
1979 1899 1978 1001
1981 1941 1979 0110
1997 1937 1979 0110
1998 x2 x1 1001
1999 x3 1998 1001
2000 1957 1999 1001
2001 1896 2000 0111
2002 1997 1999 1001
1961 1979 1981 