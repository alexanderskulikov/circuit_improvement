3 4 1
x1 x2 x3
z0 x2 x3 0110
z1 x3 z0 0111
z2 x1 z1 0100
z3 z0 z2 0110
z3