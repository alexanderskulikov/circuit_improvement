15 73 15
x1 x2 x3 x4 x5 x6 x7 x8 x9 x10 x11 x12 x13 x14 x15
z0 x4 x5 0110
z1 x6 x7 0110
z2 x8 x9 0110
z3 x10 x11 0110
z4 x12 x13 0110
z5 x14 x15 0110
z6 x1 x2 0110
z7 z6 x3 0110
z8 x1 x2 0001
z9 z6 x3 0001
z10 z8 z9 0110
z11 x4 z7 0110
z12 z0 z11 0111
z13 z0 z7 0110
z14 z12 z13 0110
z15 x6 z13 0110
z16 z13 z1 0110
z17 z15 z1 0010
z18 z12 z17 0110
z19 x8 z16 0110
z20 z2 z19 0111
z21 z2 z16 0110
z22 z20 z21 0110
z23 x10 z21 0110
z24 z21 z3 0110
z25 z23 z3 0010
z26 z20 z25 0110
z27 x12 z24 0110
z28 z4 z27 0111
z29 z4 z24 0110
z30 z28 z29 0110
z31 x14 z29 0110
z32 z29 z5 0110
z33 z31 z5 0010
z34 z28 z33 0110
z35 z14 z10 0110
z36 z18 z35 0111
z37 z18 z10 0110
z38 z36 z37 0110
z39 z22 z37 0110
z40 z37 z26 0110
z41 z39 z26 0010
z42 z36 z41 0110
z43 z40 z34 0110
z44 z30 z34 0010
z45 z40 z34 0001
z46 z44 z45 0110
z47 z46 z42 0110
z49 z46 z42 0001
a4 z43 zfcyq5 0111
a5 z47 zfcyq5 0111
a6 a4 a5 0001
a7 z32 zfcyq5 0111
a8 a6 a7 0001
a9 a4 a7 0111
a10 a5 a9 0111
a11 z43 z47 0111
a12 a8 a11 0111
a13 z32 a11 0111
a14 a5 a9 0001
a15 z32 z47 0111
a16 a8 a15 0111
a17 a12 a16 0001
a19 z47 zfcyq5 0001
a20 a13 zfcyq5 0001
a21 a11 zfcyq5 0001
a22 z32 a19 0001
a23 z43 a22 0001
a24 z43 a19 0001
a25 a15 a21 0001
a26 a22 a24 0111
zfcyq4 z42 z38 0100
zfcyq5 z49 zfcyq4 0111
a23 a24 a26 a19 a25 a21 a20 zfcyq5 a8 a6 a14 a5 a17 a12 a10