6 12 1
x1 x2 x3 x4 x5 x6 
z0 x3 x2 1001
z1 z0 x1 0111
z2 z1 x4 0110
z3 z2 x1 0110
z4 z3 x3 0110
z5 z4 z1 0001
z6 z5 x5 1001
z7 z2 z6 1001
z8 z7 z5 0010
z9 x6 z6 1011
z10 z8 x6 1001
z11 z9 z10 0001
z11 