4 8 3
x1 x2 x3 x4 
z0 x1 x3 0110
z1 x1 z0 1101
z2 x2 x4 0110
z3 z1 z2 1101
z4 x1 z3 1110
z5 z0 z2 1001
z6 x2 z5 1110
z7 z4 z6 0110
z7 z0 z3 