12 41 4
x1 x2 x3 x4 x5 x6 x7 x8 x9 x10 x11 x12
z0 x1 x2 0110
z1 z0 x3 0110
z2 x1 x2 0001
z3 z0 x3 0001
z4 z2 z3 0110
z5 x4 x5 0110
z6 x6 x7 0110
z7 x4 z1 0110
z8 z5 z7 0111
z9 z5 z1 0110
z10 z8 z9 0110
z11 x6 z9 0110
z12 z9 z6 0110
z13 z11 z6 0010
z14 z8 z13 0110
z15 x8 x9 0110
z16 x10 x11 0110
z17 x8 z12 0110
z18 z15 z17 0111
z19 z15 z12 0110
z20 z18 z19 0110
z21 x10 z19 0110
z22 z19 z16 0110
z23 z21 z16 0010
z24 z18 z23 0110
z25 z22 x12 0110
z26 z22 x12 0001
z27 z10 z4 0110
z28 z14 z27 0111
z29 z14 z4 0110
z30 z28 z29 0110
z31 z20 z29 0110
z32 z29 z24 0110
z33 z31 z24 0010
z34 z28 z33 0110
z35 z26 z32 0110
z36 z26 z32 0001
z37 z36 z34 0110
z38 z30 z34 0010
z39 z36 z34 0001
z40 z38 z39 0110
z25 z35 z37 z40