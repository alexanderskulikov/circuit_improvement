7 17 1
x1 x2 x3 x4 x5 x6 x7
z3 b6 x3 0110
b6 x2 x1 0110
z5 x4 z3 0110
z6 x4 x5 0110
z8 z3 z6 0110
z14 d5 x7 0110
a6 z3 c6 1101
c6 b7 c5 0110
a8 a6 b7 1000
b7 b5 b6 0111
b5 x3 x1 0110
a9 d8 a8 0010
c5 z5 z6 0010
d5 z8 x6 0110
d6 z8 x7 1110
d7 c6 d6 1001
d8 z14 d7 0001
a9